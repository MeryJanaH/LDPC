--**********************************************************--
-- ENSA FES --
-- Fili�re : GSEII2
--**********************************************************--
--Title : Min-Sum Algorithme
--Block : CNPU
--*************************************************************--
--File : SRC
--*************************************************************--
--                             Used Libraries
--*************************************************************--

	library ieee_proposed;
	use ieee_proposed.fixed_pkg.all;

	LIBRARY WORK;
	USE WORK.mem_types.ALL;

	
	LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;

--****************************************************--
--					ENTITY DECLARATION
--****************************************************--

ENTITY CNPU IS PORT(
	count_layer	   : IN   STD_LOGIC_VECTOR(3 DOWNTO 0);
	vnpu_out  	   : IN   T(18 DOWNTO 0);
	cnpu_out  	   : OUT  T(18 DOWNTO 0));
END CNPU;

-- **********************************************************************
-- *                        RTL Description                             *
-- **********************************************************************

ARCHITECTURE RTL OF CNPU IS 

SIGNAL mod2_in : T(15 DOWNTO 0) := (("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"));


COMPONENT mod1 IS
	PORT(
    switch_in     : IN  T(15 DOWNTO 0);
    countLayer    : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
    mod1_out      : OUT T(15 DOWNTO 0));
END COMPONENT;

COMPONENT mod2 IS
	PORT(
    mod2_in     : IN  T(18 DOWNTO 0);
    mod2_out    : OUT T(18 DOWNTO 0));
END COMPONENT;

BEGIN                 

    Md1 : mod1 PORT MAP(
	        switch_in(0)(0)   =>  vnpu_out(3)(0),
	        switch_in(1)(0)   =>  vnpu_out(4)(0),
	        switch_in(2)(0)   =>  vnpu_out(5)(0),
	        switch_in(3)(0)   =>  vnpu_out(6)(0),
	        switch_in(4)(0)   =>  vnpu_out(7)(0),
	        switch_in(5)(0)   =>  vnpu_out(8)(0),
	        switch_in(6)(0)   =>  vnpu_out(9)(0),
	        switch_in(7)(0)   =>  vnpu_out(10)(0),
	        switch_in(8)(0)   =>  vnpu_out(11)(0),
	        switch_in(9)(0)   =>  vnpu_out(12)(0),
	        switch_in(10)(0)  =>  vnpu_out(13)(0),
	        switch_in(11)(0)  =>  vnpu_out(14)(0),
	        switch_in(12)(0)  =>  vnpu_out(15)(0),
	        switch_in(13)(0)  =>  vnpu_out(16)(0),
	        switch_in(14)(0)  =>  vnpu_out(17)(0),
	        switch_in(15)(0)  =>  vnpu_out(18)(0),
	        switch_in(0)(1)   =>  vnpu_out(3)(1),
	        switch_in(1)(1)   =>  vnpu_out(4)(1),
	        switch_in(2)(1)   =>  vnpu_out(5)(1),
	        switch_in(3)(1)   =>  vnpu_out(6)(1),
	        switch_in(4)(1)   =>  vnpu_out(7)(1),
	        switch_in(5)(1)   =>  vnpu_out(8)(1),
	        switch_in(6)(1)   =>  vnpu_out(9)(1),
	        switch_in(7)(1)   =>  vnpu_out(10)(1),
	        switch_in(8)(1)   =>  vnpu_out(11)(1),
	        switch_in(9)(1)   =>  vnpu_out(12)(1),
	        switch_in(10)(1)  =>  vnpu_out(13)(1),
	        switch_in(11)(1)  =>  vnpu_out(14)(1),
	        switch_in(12)(1)  =>  vnpu_out(15)(1),
	        switch_in(13)(1)  =>  vnpu_out(16)(1),
	        switch_in(14)(1)  =>  vnpu_out(17)(1),
	        switch_in(15)(1)  =>  vnpu_out(18)(1),
	        switch_in(0)(2)   =>  vnpu_out(3)(2),
	        switch_in(1)(2)   =>  vnpu_out(4)(2),
	        switch_in(2)(2)   =>  vnpu_out(5)(2),
	        switch_in(3)(2)   =>  vnpu_out(6)(2),
	        switch_in(4)(2)   =>  vnpu_out(7)(2),
	        switch_in(5)(2)   =>  vnpu_out(8)(2),
	        switch_in(6)(2)   =>  vnpu_out(9)(2),
	        switch_in(7)(2)   =>  vnpu_out(10)(2),
	        switch_in(8)(2)   =>  vnpu_out(11)(2),
	        switch_in(9)(2)   =>  vnpu_out(12)(2),
	        switch_in(10)(2)  =>  vnpu_out(13)(2),
	        switch_in(11)(2)  =>  vnpu_out(14)(2),
	        switch_in(12)(2)  =>  vnpu_out(15)(2),
	        switch_in(13)(2)  =>  vnpu_out(16)(2),
	        switch_in(14)(2)  =>  vnpu_out(17)(2),
	        switch_in(15)(2)  =>  vnpu_out(18)(2),
	        switch_in(0)(3)   =>  vnpu_out(3)(3),
	        switch_in(1)(3)   =>  vnpu_out(4)(3),
	        switch_in(2)(3)   =>  vnpu_out(5)(3),
	        switch_in(3)(3)   =>  vnpu_out(6)(3),
	        switch_in(4)(3)   =>  vnpu_out(7)(3),
	        switch_in(5)(3)   =>  vnpu_out(8)(3),
	        switch_in(6)(3)   =>  vnpu_out(9)(3),
	        switch_in(7)(3)   =>  vnpu_out(10)(3),
	        switch_in(8)(3)   =>  vnpu_out(11)(3),
	        switch_in(9)(3)   =>  vnpu_out(12)(3),
	        switch_in(10)(3)  =>  vnpu_out(13)(3),
	        switch_in(11)(3)  =>  vnpu_out(14)(3),
	        switch_in(12)(3)  =>  vnpu_out(15)(3),
	        switch_in(13)(3)  =>  vnpu_out(16)(3),
	        switch_in(14)(3)  =>  vnpu_out(17)(3),
	        switch_in(15)(3)  =>  vnpu_out(18)(3),
	        switch_in(0)(4)   =>  vnpu_out(3)(4),
	        switch_in(1)(4)   =>  vnpu_out(4)(4),
	        switch_in(2)(4)   =>  vnpu_out(5)(4),
	        switch_in(3)(4)   =>  vnpu_out(6)(4),
	        switch_in(4)(4)   =>  vnpu_out(7)(4),
	        switch_in(5)(4)   =>  vnpu_out(8)(4),
	        switch_in(6)(4)   =>  vnpu_out(9)(4),
	        switch_in(7)(4)   =>  vnpu_out(10)(4),
	        switch_in(8)(4)   =>  vnpu_out(11)(4),
	        switch_in(9)(4)   =>  vnpu_out(12)(4),
	        switch_in(10)(4)  =>  vnpu_out(13)(4),
	        switch_in(11)(4)  =>  vnpu_out(14)(4),
	        switch_in(12)(4)  =>  vnpu_out(15)(4),
	        switch_in(13)(4)  =>  vnpu_out(16)(4),
	        switch_in(14)(4)  =>  vnpu_out(17)(4),
	        switch_in(15)(4)  =>  vnpu_out(18)(4),
	        switch_in(0)(5)   =>  vnpu_out(3)(5),
	        switch_in(1)(5)   =>  vnpu_out(4)(5),
	        switch_in(2)(5)   =>  vnpu_out(5)(5),
	        switch_in(3)(5)   =>  vnpu_out(6)(5),
	        switch_in(4)(5)   =>  vnpu_out(7)(5),
	        switch_in(5)(5)   =>  vnpu_out(8)(5),
	        switch_in(6)(5)   =>  vnpu_out(9)(5),
	        switch_in(7)(5)   =>  vnpu_out(10)(5),
	        switch_in(8)(5)   =>  vnpu_out(11)(5),
	        switch_in(9)(5)   =>  vnpu_out(12)(5),
	        switch_in(10)(5)  =>  vnpu_out(13)(5),
	        switch_in(11)(5)  =>  vnpu_out(14)(5),
	        switch_in(12)(5)  =>  vnpu_out(15)(5),
	        switch_in(13)(5)  =>  vnpu_out(16)(5),
	        switch_in(14)(5)  =>  vnpu_out(17)(5),
	        switch_in(15)(5)  =>  vnpu_out(18)(5),
	        switch_in(0)(6)   =>  vnpu_out(3)(6),
	        switch_in(1)(6)   =>  vnpu_out(4)(6),
	        switch_in(2)(6)   =>  vnpu_out(5)(6),
	        switch_in(3)(6)   =>  vnpu_out(6)(6),
	        switch_in(4)(6)   =>  vnpu_out(7)(6),
	        switch_in(5)(6)   =>  vnpu_out(8)(6),
	        switch_in(6)(6)   =>  vnpu_out(9)(6),
	        switch_in(7)(6)   =>  vnpu_out(10)(6),
	        switch_in(8)(6)   =>  vnpu_out(11)(6),
	        switch_in(9)(6)   =>  vnpu_out(12)(6),
	        switch_in(10)(6)  =>  vnpu_out(13)(6),
	        switch_in(11)(6)  =>  vnpu_out(14)(6),
	        switch_in(12)(6)  =>  vnpu_out(15)(6),
	        switch_in(13)(6)  =>  vnpu_out(16)(6),
	        switch_in(14)(6)  =>  vnpu_out(17)(6),
	        switch_in(15)(6)  =>  vnpu_out(18)(6),
	        switch_in(0)(7)   =>  vnpu_out(3)(7),
	        switch_in(1)(7)   =>  vnpu_out(4)(7),
	        switch_in(2)(7)   =>  vnpu_out(5)(7),
	        switch_in(3)(7)   =>  vnpu_out(6)(7),
	        switch_in(4)(7)   =>  vnpu_out(7)(7),
	        switch_in(5)(7)   =>  vnpu_out(8)(7),
	        switch_in(6)(7)   =>  vnpu_out(9)(7),
	        switch_in(7)(7)   =>  vnpu_out(10)(7),
	        switch_in(8)(7)   =>  vnpu_out(11)(7),
	        switch_in(9)(7)   =>  vnpu_out(12)(7),
	        switch_in(10)(7)  =>  vnpu_out(13)(7),
	        switch_in(11)(7)  =>  vnpu_out(14)(7),
	        switch_in(12)(7)  =>  vnpu_out(15)(7),
	        switch_in(13)(7)  =>  vnpu_out(16)(7),
	        switch_in(14)(7)  =>  vnpu_out(17)(7),
	        switch_in(15)(7)  =>  vnpu_out(18)(7),
            countLayer  	  => count_layer,
	        mod1_out(0)(0)   =>  mod2_in(0)(0),
	        mod1_out(1)(0)   =>  mod2_in(1)(0),
	        mod1_out(2)(0)   =>  mod2_in(2)(0),
	        mod1_out(3)(0)   =>  mod2_in(3)(0),
	        mod1_out(4)(0)   =>  mod2_in(4)(0),
	        mod1_out(5)(0)   =>  mod2_in(5)(0),
	        mod1_out(6)(0)   =>  mod2_in(6)(0),
	        mod1_out(7)(0)   =>  mod2_in(7)(0),
	        mod1_out(8)(0)   =>  mod2_in(8)(0),
	        mod1_out(9)(0)   =>  mod2_in(9)(0),
	        mod1_out(10)(0)  =>  mod2_in(10)(0),
	        mod1_out(11)(0)  =>  mod2_in(11)(0),
	        mod1_out(12)(0)  =>  mod2_in(12)(0),
	        mod1_out(13)(0)  =>  mod2_in(13)(0),
	        mod1_out(14)(0)  =>  mod2_in(14)(0),
	        mod1_out(15)(0)  =>  mod2_in(15)(0),
	        mod1_out(0)(1)   =>  mod2_in(0)(1),
	        mod1_out(1)(1)   =>  mod2_in(1)(1),
	        mod1_out(2)(1)   =>  mod2_in(2)(1),
	        mod1_out(3)(1)   =>  mod2_in(3)(1),
	        mod1_out(4)(1)   =>  mod2_in(4)(1),
	        mod1_out(5)(1)   =>  mod2_in(5)(1),
	        mod1_out(6)(1)   =>  mod2_in(6)(1),
	        mod1_out(7)(1)   =>  mod2_in(7)(1),
	        mod1_out(8)(1)   =>  mod2_in(8)(1),
	        mod1_out(9)(1)   =>  mod2_in(9)(1),
	        mod1_out(10)(1)  =>  mod2_in(10)(1),
	        mod1_out(11)(1)  =>  mod2_in(11)(1),
	        mod1_out(12)(1)  =>  mod2_in(12)(1),
	        mod1_out(13)(1)  =>  mod2_in(13)(1),
	        mod1_out(14)(1)  =>  mod2_in(14)(1),
	        mod1_out(15)(1)  =>  mod2_in(15)(1),
	        mod1_out(0)(2)   =>  mod2_in(0)(2),
	        mod1_out(1)(2)   =>  mod2_in(1)(2),
	        mod1_out(2)(2)   =>  mod2_in(2)(2),
	        mod1_out(3)(2)   =>  mod2_in(3)(2),
	        mod1_out(4)(2)   =>  mod2_in(4)(2),
	        mod1_out(5)(2)   =>  mod2_in(5)(2),
	        mod1_out(6)(2)   =>  mod2_in(6)(2),
	        mod1_out(7)(2)   =>  mod2_in(7)(2),
	        mod1_out(8)(2)   =>  mod2_in(8)(2),
	        mod1_out(9)(2)   =>  mod2_in(9)(2),
	        mod1_out(10)(2)  =>  mod2_in(10)(2),
	        mod1_out(11)(2)  =>  mod2_in(11)(2),
	        mod1_out(12)(2)  =>  mod2_in(12)(2),
	        mod1_out(13)(2)  =>  mod2_in(13)(2),
	        mod1_out(14)(2)  =>  mod2_in(14)(2),
	        mod1_out(15)(2)  =>  mod2_in(15)(2),
	        mod1_out(0)(3)   =>  mod2_in(0)(3),
	        mod1_out(1)(3)   =>  mod2_in(1)(3),
	        mod1_out(2)(3)   =>  mod2_in(2)(3),
	        mod1_out(3)(3)   =>  mod2_in(3)(3),
	        mod1_out(4)(3)   =>  mod2_in(4)(3),
	        mod1_out(5)(3)   =>  mod2_in(5)(3),
	        mod1_out(6)(3)   =>  mod2_in(6)(3),
	        mod1_out(7)(3)   =>  mod2_in(7)(3),
	        mod1_out(8)(3)   =>  mod2_in(8)(3),
	        mod1_out(9)(3)   =>  mod2_in(9)(3),
	        mod1_out(10)(3)  =>  mod2_in(10)(3),
	        mod1_out(11)(3)  =>  mod2_in(11)(3),
	        mod1_out(12)(3)  =>  mod2_in(12)(3),
	        mod1_out(13)(3)  =>  mod2_in(13)(3),
	        mod1_out(14)(3)  =>  mod2_in(14)(3),
	        mod1_out(15)(3)  =>  mod2_in(15)(3),
	        mod1_out(0)(4)   =>  mod2_in(0)(4),
	        mod1_out(1)(4)   =>  mod2_in(1)(4),
	        mod1_out(2)(4)   =>  mod2_in(2)(4),
	        mod1_out(3)(4)   =>  mod2_in(3)(4),
	        mod1_out(4)(4)   =>  mod2_in(4)(4),
	        mod1_out(5)(4)   =>  mod2_in(5)(4),
	        mod1_out(6)(4)   =>  mod2_in(6)(4),
	        mod1_out(7)(4)   =>  mod2_in(7)(4),
	        mod1_out(8)(4)   =>  mod2_in(8)(4),
	        mod1_out(9)(4)   =>  mod2_in(9)(4),
	        mod1_out(10)(4)  =>  mod2_in(10)(4),
	        mod1_out(11)(4)  =>  mod2_in(11)(4),
	        mod1_out(12)(4)  =>  mod2_in(12)(4),
	        mod1_out(13)(4)  =>  mod2_in(13)(4),
	        mod1_out(14)(4)  =>  mod2_in(14)(4),
	        mod1_out(15)(4)  =>  mod2_in(15)(4),
	        mod1_out(0)(5)   =>  mod2_in(0)(5),
	        mod1_out(1)(5)   =>  mod2_in(1)(5),
	        mod1_out(2)(5)   =>  mod2_in(2)(5),
	        mod1_out(3)(5)   =>  mod2_in(3)(5),
	        mod1_out(4)(5)   =>  mod2_in(4)(5),
	        mod1_out(5)(5)   =>  mod2_in(5)(5),
	        mod1_out(6)(5)   =>  mod2_in(6)(5),
	        mod1_out(7)(5)   =>  mod2_in(7)(5),
	        mod1_out(8)(5)   =>  mod2_in(8)(5),
	        mod1_out(9)(5)   =>  mod2_in(9)(5),
	        mod1_out(10)(5)  =>  mod2_in(10)(5),
	        mod1_out(11)(5)  =>  mod2_in(11)(5),
	        mod1_out(12)(5)  =>  mod2_in(12)(5),
	        mod1_out(13)(5)  =>  mod2_in(13)(5),
	        mod1_out(14)(5)  =>  mod2_in(14)(5),
	        mod1_out(15)(5)  =>  mod2_in(15)(5),
	        mod1_out(0)(6)   =>  mod2_in(0)(6),
	        mod1_out(1)(6)   =>  mod2_in(1)(6),
	        mod1_out(2)(6)   =>  mod2_in(2)(6),
	        mod1_out(3)(6)   =>  mod2_in(3)(6),
	        mod1_out(4)(6)   =>  mod2_in(4)(6),
	        mod1_out(5)(6)   =>  mod2_in(5)(6),
	        mod1_out(6)(6)   =>  mod2_in(6)(6),
	        mod1_out(7)(6)   =>  mod2_in(7)(6),
	        mod1_out(8)(6)   =>  mod2_in(8)(6),
	        mod1_out(9)(6)   =>  mod2_in(9)(6),
	        mod1_out(10)(6)  =>  mod2_in(10)(6),
	        mod1_out(11)(6)  =>  mod2_in(11)(6),
	        mod1_out(12)(6)  =>  mod2_in(12)(6),
	        mod1_out(13)(6)  =>  mod2_in(13)(6),
	        mod1_out(14)(6)  =>  mod2_in(14)(6),
	        mod1_out(15)(6)  =>  mod2_in(15)(6),
	        mod1_out(0)(7)   =>  mod2_in(0)(7),
	        mod1_out(1)(7)   =>  mod2_in(1)(7),
	        mod1_out(2)(7)   =>  mod2_in(2)(7),
	        mod1_out(3)(7)   =>  mod2_in(3)(7),
	        mod1_out(4)(7)   =>  mod2_in(4)(7),
	        mod1_out(5)(7)   =>  mod2_in(5)(7),
	        mod1_out(6)(7)   =>  mod2_in(6)(7),
	        mod1_out(7)(7)   =>  mod2_in(7)(7),
	        mod1_out(8)(7)   =>  mod2_in(8)(7),
	        mod1_out(9)(7)   =>  mod2_in(9)(7),
	        mod1_out(10)(7)  =>  mod2_in(10)(7),
	        mod1_out(11)(7)  =>  mod2_in(11)(7),
	        mod1_out(12)(7)  =>  mod2_in(12)(7),
	        mod1_out(13)(7)  =>  mod2_in(13)(7),
	        mod1_out(14)(7)  =>  mod2_in(14)(7),
	        mod1_out(15)(7)  =>  mod2_in(15)(7));
  
    Md2 : mod2 PORT MAP(
            mod2_in(0)(0)   =>  vnpu_out(0)(0),
	        mod2_in(1)(0)   =>  vnpu_out(1)(0),
	        mod2_in(2)(0)   =>  vnpu_out(2)(0),
	        mod2_in(3)(0)   =>  mod2_in(0)(0),
	        mod2_in(4)(0)   =>  mod2_in(1)(0),
	        mod2_in(5)(0)   =>  mod2_in(2)(0),
	        mod2_in(6)(0)   =>  mod2_in(3)(0),
	        mod2_in(7)(0)   =>  mod2_in(4)(0),
	        mod2_in(8)(0)   =>  mod2_in(5)(0),
	        mod2_in(9)(0)   =>  mod2_in(6)(0),
	        mod2_in(10)(0)  =>  mod2_in(7)(0),
	        mod2_in(11)(0)  =>  mod2_in(8)(0),
	        mod2_in(12)(0)  =>  mod2_in(9)(0),
	        mod2_in(13)(0)  =>  mod2_in(10)(0),
	        mod2_in(14)(0)  =>  mod2_in(11)(0),
	        mod2_in(15)(0)  =>  mod2_in(12)(0),
	        mod2_in(16)(0)  =>  mod2_in(13)(0),
	        mod2_in(17)(0)  =>  mod2_in(14)(0),
	        mod2_in(18)(0)  =>  mod2_in(15)(0),
	        mod2_in(0)(1)   =>  vnpu_out(0)(1),
	        mod2_in(1)(1)   =>  vnpu_out(1)(1),
	        mod2_in(2)(1)   =>  vnpu_out(2)(1),
	        mod2_in(3)(1)   =>  mod2_in(0)(1),
	        mod2_in(4)(1)   =>  mod2_in(1)(1),
	        mod2_in(5)(1)   =>  mod2_in(2)(1),
	        mod2_in(6)(1)   =>  mod2_in(3)(1),
	        mod2_in(7)(1)   =>  mod2_in(4)(1),
	        mod2_in(8)(1)   =>  mod2_in(5)(1),
	        mod2_in(9)(1)   =>  mod2_in(6)(1),
	        mod2_in(10)(1)  =>  mod2_in(7)(1),
	        mod2_in(11)(1)  =>  mod2_in(8)(1),
	        mod2_in(12)(1)  =>  mod2_in(9)(1),
	        mod2_in(13)(1)  =>  mod2_in(10)(1),
	        mod2_in(14)(1)  =>  mod2_in(11)(1),
	        mod2_in(15)(1)  =>  mod2_in(12)(1),
	        mod2_in(16)(1)  =>  mod2_in(13)(1),
	        mod2_in(17)(1)  =>  mod2_in(14)(1),
	        mod2_in(18)(1)  =>  mod2_in(15)(1),
	        mod2_in(0)(2)   =>  vnpu_out(0)(2),
	        mod2_in(1)(2)   =>  vnpu_out(1)(2),
	        mod2_in(2)(2)   =>  vnpu_out(2)(2),
	        mod2_in(3)(2)   =>  mod2_in(0)(2),
	        mod2_in(4)(2)   =>  mod2_in(1)(2),
	        mod2_in(5)(2)   =>  mod2_in(2)(2),
	        mod2_in(6)(2)   =>  mod2_in(3)(2),
	        mod2_in(7)(2)   =>  mod2_in(4)(2),
	        mod2_in(8)(2)   =>  mod2_in(5)(2),
	        mod2_in(9)(2)   =>  mod2_in(6)(2),
	        mod2_in(10)(2)  =>  mod2_in(7)(2),
	        mod2_in(11)(2)  =>  mod2_in(8)(2),
	        mod2_in(12)(2)  =>  mod2_in(9)(2),
	        mod2_in(13)(2)  =>  mod2_in(10)(2),
	        mod2_in(14)(2)  =>  mod2_in(11)(2),
	        mod2_in(15)(2)  =>  mod2_in(12)(2),
	        mod2_in(16)(2)  =>  mod2_in(13)(2),
	        mod2_in(17)(2)  =>  mod2_in(14)(2),
	        mod2_in(18)(2)  =>  mod2_in(15)(2),
	        mod2_in(0)(3)   =>  vnpu_out(0)(3),
	        mod2_in(1)(3)   =>  vnpu_out(1)(3),
	        mod2_in(2)(3)   =>  vnpu_out(2)(3),
	        mod2_in(3)(3)   =>  mod2_in(0)(3),
	        mod2_in(4)(3)   =>  mod2_in(1)(3),
	        mod2_in(5)(3)   =>  mod2_in(2)(3),
	        mod2_in(6)(3)   =>  mod2_in(3)(3),
	        mod2_in(7)(3)   =>  mod2_in(4)(3),
	        mod2_in(8)(3)   =>  mod2_in(5)(3),
	        mod2_in(9)(3)   =>  mod2_in(6)(3),
	        mod2_in(10)(3)  =>  mod2_in(7)(3),
	        mod2_in(11)(3)  =>  mod2_in(8)(3),
	        mod2_in(12)(3)  =>  mod2_in(9)(3),
	        mod2_in(13)(3)  =>  mod2_in(10)(3),
	        mod2_in(14)(3)  =>  mod2_in(11)(3),
	        mod2_in(15)(3)  =>  mod2_in(12)(3),
	        mod2_in(16)(3)  =>  mod2_in(13)(3),
	        mod2_in(17)(3)  =>  mod2_in(14)(3),
	        mod2_in(18)(3)  =>  mod2_in(15)(3),
	        mod2_in(0)(4)   =>  vnpu_out(0)(4),
	        mod2_in(1)(4)   =>  vnpu_out(1)(4),
	        mod2_in(2)(4)   =>  vnpu_out(2)(4),
	        mod2_in(3)(4)   =>  mod2_in(0)(4),
	        mod2_in(4)(4)   =>  mod2_in(1)(4),
	        mod2_in(5)(4)   =>  mod2_in(2)(4),
	        mod2_in(6)(4)   =>  mod2_in(3)(4),
	        mod2_in(7)(4)   =>  mod2_in(4)(4),
	        mod2_in(8)(4)   =>  mod2_in(5)(4),
	        mod2_in(9)(4)   =>  mod2_in(6)(4),
	        mod2_in(10)(4)  =>  mod2_in(7)(4),
	        mod2_in(11)(4)  =>  mod2_in(8)(4),
	        mod2_in(12)(4)  =>  mod2_in(9)(4),
	        mod2_in(13)(4)  =>  mod2_in(10)(4),
	        mod2_in(14)(4)  =>  mod2_in(11)(4),
	        mod2_in(15)(4)  =>  mod2_in(12)(4),
	        mod2_in(16)(4)  =>  mod2_in(13)(4),
	        mod2_in(17)(4)  =>  mod2_in(14)(4),
	        mod2_in(18)(4)  =>  mod2_in(15)(4),
	        mod2_in(0)(5)   =>  vnpu_out(0)(5),
	        mod2_in(1)(5)   =>  vnpu_out(1)(5),
	        mod2_in(2)(5)   =>  vnpu_out(2)(5),
	        mod2_in(3)(5)   =>  mod2_in(0)(5),
	        mod2_in(4)(5)   =>  mod2_in(1)(5),
	        mod2_in(5)(5)   =>  mod2_in(2)(5),
	        mod2_in(6)(5)   =>  mod2_in(3)(5),
	        mod2_in(7)(5)   =>  mod2_in(4)(5),
	        mod2_in(8)(5)   =>  mod2_in(5)(5),
	        mod2_in(9)(5)   =>  mod2_in(6)(5),
	        mod2_in(10)(5)  =>  mod2_in(7)(5),
	        mod2_in(11)(5)  =>  mod2_in(8)(5),
	        mod2_in(12)(5)  =>  mod2_in(9)(5),
	        mod2_in(13)(5)  =>  mod2_in(10)(5),
	        mod2_in(14)(5)  =>  mod2_in(11)(5),
	        mod2_in(15)(5)  =>  mod2_in(12)(5),
	        mod2_in(16)(5)  =>  mod2_in(13)(5),
	        mod2_in(17)(5)  =>  mod2_in(14)(5),
	        mod2_in(18)(5)  =>  mod2_in(15)(5),
	        mod2_in(0)(6)   =>  vnpu_out(0)(6),
	        mod2_in(1)(6)   =>  vnpu_out(1)(6),
	        mod2_in(2)(6)   =>  vnpu_out(2)(6),
	        mod2_in(3)(6)   =>  mod2_in(0)(6),
	        mod2_in(4)(6)   =>  mod2_in(1)(6),
	        mod2_in(5)(6)   =>  mod2_in(2)(6),
	        mod2_in(6)(6)   =>  mod2_in(3)(6),
	        mod2_in(7)(6)   =>  mod2_in(4)(6),
	        mod2_in(8)(6)   =>  mod2_in(5)(6),
	        mod2_in(9)(6)   =>  mod2_in(6)(6),
	        mod2_in(10)(6)  =>  mod2_in(7)(6),
	        mod2_in(11)(6)  =>  mod2_in(8)(6),
	        mod2_in(12)(6)  =>  mod2_in(9)(6),
	        mod2_in(13)(6)  =>  mod2_in(10)(6),
	        mod2_in(14)(6)  =>  mod2_in(11)(6),
	        mod2_in(15)(6)  =>  mod2_in(12)(6),
	        mod2_in(16)(6)  =>  mod2_in(13)(6),
	        mod2_in(17)(6)  =>  mod2_in(14)(6),
	        mod2_in(18)(6)  =>  mod2_in(15)(6),
	        mod2_in(0)(7)   =>  vnpu_out(0)(7),
	        mod2_in(1)(7)   =>  vnpu_out(1)(7),
	        mod2_in(2)(7)   =>  vnpu_out(2)(7),
	        mod2_in(3)(7)   =>  mod2_in(0)(7),
	        mod2_in(4)(7)   =>  mod2_in(1)(7),
	        mod2_in(5)(7)   =>  mod2_in(2)(7),
	        mod2_in(6)(7)   =>  mod2_in(3)(7),
	        mod2_in(7)(7)   =>  mod2_in(4)(7),
	        mod2_in(8)(7)   =>  mod2_in(5)(7),
	        mod2_in(9)(7)   =>  mod2_in(6)(7),
	        mod2_in(10)(7)  =>  mod2_in(7)(7),
	        mod2_in(11)(7)  =>  mod2_in(8)(7),
	        mod2_in(12)(7)  =>  mod2_in(9)(7),
	        mod2_in(13)(7)  =>  mod2_in(10)(7),
	        mod2_in(14)(7)  =>  mod2_in(11)(7),
	        mod2_in(15)(7)  =>  mod2_in(12)(7),
	        mod2_in(16)(7)  =>  mod2_in(13)(7),
	        mod2_in(17)(7)  =>  mod2_in(14)(7),
	        mod2_in(18)(7)  =>  mod2_in(15)(7),
            mod2_out        => cnpu_out);
                     
END RTL;
