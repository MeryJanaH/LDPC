--***********************************************************************************************************--
--						USED LIBRAIRIES						     --
--***********************************************************************************************************--
LIBRARY ieee_proposed;
USE ieee_proposed.fixed_pkg.all;
USE WORK.mem_types.ALL;
--*****************************************************************************************************************--
--						ENTITY DECLARATION						   --
--*****************************************************************************************************************--
ENTITY conv_T2Tb IS PORT(
	R: IN T(18 DOWNTO 0);
	S : OUT Tb(18 DOWNTO 0)
);
END conv_T2Tb;
--*****************************************************************************************************************--
--						ARCHITECTURE DESCRIPTION					   --
--*****************************************************************************************************************--
ARCHITECTURE RTL OF conv_T2Tb IS
BEGIN
	PROCESS(R)
	BEGIN
		FOR i IN 18 DOWNTO 0 LOOP
			FOR j IN 7 DOWNTO 0 LOOP
				S(i)(j) <= resize(R(i)(j),3,-7);
			END LOOP;
		END LOOP;
	END PROCESS;
END RTL;