--***********************************************************************************************************--
--						USED LIBRAIRIES						     --
--***********************************************************************************************************--
USE WORK.mem_types.ALL;
--**********************************************************************************************************--
--						ENTITY DECLARATION					    --
--**********************************************************************************************************--
ENTITY inter_wt_19 IS
PORT( 
	N: IN T(18 DOWNTO 0);
	R: IN T(15 DOWNTO 0);
	Ind: IN index(18 DOWNTO 0);
	S: OUT T(34 DOWNTO 0)
);
END inter_wt_19;
--***********************************************************************************************************--
--						ARCHITECTURE DESCRIPTION				     --
--***********************************************************************************************************--
ARCHITECTURE RTL OF inter_wt_19 IS
BEGIN
	PROCESS(N,R)
	VARIABLE j : INTEGER;
	VARIABLE k : INTEGER;
	BEGIN
		j:=18;
		k:=15;
		FOR i IN 34 DOWNTO 0 LOOP
			IF  j>=0 and Ind(j)=i THEN
				S(i)<= N(j);
				j:=j-1;
			ELSIF  k>=0 THEN
				S(i)<= R(k) ;
				k:=k-1;
			END IF;
		END LOOP;
	END PROCESS;
END RTL;
	 