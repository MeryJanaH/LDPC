--***********************************************************************************************************--
--						USED LIBRAIRIES						     --
--***********************************************************************************************************--
USE WORK.mem_types.ALL;
--**********************************************************************************************************--
--						ENTITY DECLARATION					    --
--**********************************************************************************************************--
ENTITY up_down IS PORT(
	A: IN T(18 DOWNTO 0);
	S: OUT T(18 DOWNTO 0));
END up_down;
--***********************************************************************************************************--
--						ARCHITECTURE DESCRIPTION				     --
--***********************************************************************************************************--
ARCHITECTURE RTL OF up_down IS
BEGIN
	PROCESS(A)
	VARIABLE j: INTEGER;
	BEGIN
		j:=0;
		FOR i IN 18 DOWNTO 0 LOOP
			S(j)<= A(i);
			j:=j+1;
		END LOOP;		
	END PROCESS;
END RTL;