--*****************************************************************************************************************--
--						USED LIBRAIRIES							   --
--*****************************************************************************************************************--
USE WORK.mem_types.ALL;
--*****************************************************************************************************************--
--						ENTITY DECLARATION						   --
--*****************************************************************************************************************--
ENTITY control_filter_19 IS PORT(
	C: IN control;
	S: OUT shift);
END control_filter_19;
--*****************************************************************************************************************--
--						ARCHITECTURE DESCRIPTION					   --
--*****************************************************************************************************************--
ARCHITECTURE RTL OF control_filter_19 IS
BEGIN
	PROCESS(C)
	VARIABLE j: integer;
	BEGIN
		j:=18;
		FOR i IN 34 DOWNTO 0 LOOP
			IF C(i) >= 0 THEN
					S(j)<= C(i);
					j:=j-1;
			END IF;
		END LOOP;
		WHILE j>-1 LOOP
			S(j)<= 0;
			j:=j-1;
		END LOOP;
	END PROCESS;
END RTL ;