--***********************************************************************************************************--
--						USED LIBRAIRIES						     --
--***********************************************************************************************************--
USE WORK.mem_types.ALL;
--**********************************************************************************************************--
--						ENTITY DECLARATION					    --
--**********************************************************************************************************--
ENTITY down_up IS PORT(
	A: IN T(18 DOWNTO 0);
	S: OUT T(18 DOWNTO 0));
END down_up;
--***********************************************************************************************************--
--						ARCHITECTURE DESCRIPTION				     --
--***********************************************************************************************************--
ARCHITECTURE RTL OF down_up IS
BEGIN
	PROCESS(A)
	VARIABLE j: INTEGER;
	BEGIN
		j:=0;
		FOR i IN 18 DOWNTO 0 LOOP
			S(i)<= A(j);
			j:=j+1;
		END LOOP;		
	END PROCESS;
END RTL;