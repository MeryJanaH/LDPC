--**********************************************************--
-- ENSA FES --
-- Fili�re : GSEII2
--**********************************************************--
--Title : Min-Sum Algorithme
--Block : C.G.memory 
--*************************************************************--
--*************************************************************--
--File : src
--*************************************************************--
--                             Used Libraries
--*************************************************************--

	LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
	USE IEEE.numeric_std.ALL;
	use IEEE.std_logic_unsigned.all;

	LIBRARY WORK;
	USE WORK.mem_types.ALL;
	
--************************************************************--
--                            ENTITY Declaration
--************************************************************--

ENTITY Code_gen IS PORT(  
    countLayer      : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
    mem_in  	 : IN  T(34 DOWNTO 0);
    MemAdr   	 : IN  STD_LOGIC;
    recv_LLR     : IN  T(34 DOWNTO 0);
    clk          : IN  STD_LOGIC;
	reset        : IN  STD_LOGIC;
	recv_LLR2    : OUT T(34 DOWNTO 0));  
END Code_gen;

--**********************************************************************************--
--                              RTL DESCRIPTION                                     --
--**********************************************************************************--
ARCHITECTURE RTL OF Code_gen IS
	
SIGNAL mem_o : T(34 DOWNTO 0) := (("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
			            			("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"));

COMPONENT Layer_mem IS
	PORT(
    countLayer      : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
    mem_in  	: IN   T(34 DOWNTO 0);
    mem_out   	: OUT  T(34 DOWNTO 0);
	MemAdr		: IN   STD_LOGIC;
    clk         : IN   STD_LOGIC;
	reset       : IN   STD_LOGIC);
END COMPONENT;

COMPONENT switch_mem IS
	PORT(
    recv_LLR  	 : IN  T(34 DOWNTO 0);
    Code_gen   	 : IN  T(34 DOWNTO 0);
    MemAdr		 : IN  STD_LOGIC;
    switch_out   : OUT T(34 DOWNTO 0));  
END COMPONENT;
		
BEGIN 

n1 : Layer_mem PORT MAP(
         countLayer     => countLayer,
         mem_in  => mem_in,
         mem_out => mem_o,
		 MemAdr     => MemAdr,
         clk     => clk,
         reset   => reset);
 
n2 : switch_mem PORT MAP(
         recv_LLR   => recv_LLR,
         Code_gen   => mem_o,
         MemAdr     => MemAdr,
         switch_out => recv_LLR2);
                     
END RTL;
